`timescale 1ns / 1ns

module RandomGen(Clk, Rst, RandomValue);

   input Clk, Rst;
   output [ ] RandomValue; // you need decide the number of bits here.
   
   
endmodule
